// ------------------------------------------------------------------------- --
// Title         : DCF77-Decoder
// Project       : Praktikum FPGA-Entwurfstechnik
// ------------------------------------------------------------------------- --
// File          : timeAndDateClock.v
// Author        : Tim Stadtmann
// Company       : IDS RWTH Aachen 
// Created       : 2018/09/20
// ------------------------------------------------------------------------- --
// Description   : Decodes the dcf77 signal
// ------------------------------------------------------------------------- --
// Revisions     :
// Date        Version  Author  Description
// 2018/09/20  1.0      TS      Created
// ------------------------------------------------------------------------- --

module dcf77_decoder(clk,             // Global 10MHz clock 
                     clk_en_1hz,      // Indicates start of second
                     nReset,          // Global reset
                     minute_start_in, // New minute trigger
                     dcf_Signal_in,   // DFC Signal
                     timeAndDate_out,
                     data_valid,      // Control signal, High if data is valid
                     dcf_value);      // Decoded value of dcf input signal
                     
input clk, 
      clk_en_1hz,     
      nReset,  
      minute_start_in,
      dcf_Signal_in;  
      
output reg[43:0]  timeAndDate_out;
output reg        data_valid;
output reg           dcf_value;
   
// ---------- YOUR CODE HERE ---------- 
reg minute_start_observed = 0;
reg [7:0] counter = 0;
reg [59:0]full_dcf_signal =0;
initial data_valid = 0;

reg error_1 = 1;
reg error_2 = 1;
reg error_3 = 1;


always @(posedge minute_start_in, negedge clk_en_1hz, negedge nReset) begin
	if(!nReset) begin
		counter <= 0;
		data_valid <= 0;
		full_dcf_signal <= 0;
		minute_start_observed <= 0;
	end
	else begin
	if(minute_start_in) begin
		minute_start_observed <= 1;
		full_dcf_signal[59] <= 0;
		counter <= 59;
	end
	else if(!clk_en_1hz) begin
		if(minute_start_observed) begin
			minute_start_observed <= 0;
			if(!error_1 & !error_2 & !error_3) begin
				data_valid <= 1;
			end
			counter <= 0;
			dcf_value <= ~dcf_Signal_in;
			full_dcf_signal[0] <= 0;
		end
		else begin
			data_valid <= 0;
			dcf_value <= ~dcf_Signal_in;
			counter <= counter + 1;
			full_dcf_signal[counter+1] <= ~dcf_Signal_in;
		end
	end
	end
end

always @( posedge clk, negedge nReset) begin
	if(!nReset) begin
		error_1 <= 1;
		error_2 <= 1;
		error_3 <= 1;
		timeAndDate_out <= 0;
	end
	else begin
		timeAndDate_out[13:7] <= full_dcf_signal[27:21];
		// assign hours
		timeAndDate_out[19:14] <= full_dcf_signal[34:29];
		// assign days
		timeAndDate_out[25:20]	<= full_dcf_signal[41:36];
		//weekday
		timeAndDate_out[41:39]	<= full_dcf_signal[44:42];
		//month
		timeAndDate_out[30:26]	<= full_dcf_signal[49:45];
		//year
		timeAndDate_out[38:31]	<= full_dcf_signal[57:50];
		//timezone
		timeAndDate_out[43:42] <= full_dcf_signal[18:17];
		
		if(counter[7:0] == 1) begin
			error_1 <= 1;
			error_2 <= 1;
			error_3 <= 1;
		end
		else if(counter[7:0] == 28) begin
			error_1 <= ^ full_dcf_signal[28:21];
		end
		else if(counter[7:0] == 35) begin	
			error_2 <= ^ full_dcf_signal[35:29];
		end
		else if(counter[7:0] == 58) begin
			error_3 <= ^ full_dcf_signal[58:36];
		end
	end
end
            
endmodule             
              

